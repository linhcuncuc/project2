library verilog;
use verilog.vl_types.all;
entity tb_counter1 is
end tb_counter1;
